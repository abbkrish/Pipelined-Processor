library verilog;
use verilog.vl_types.all;
entity icache_datapath_sv_unit is
end icache_datapath_sv_unit;
