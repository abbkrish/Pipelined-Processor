library verilog;
use verilog.vl_types.all;
entity MP3_sv_unit is
end MP3_sv_unit;
