library verilog;
use verilog.vl_types.all;
entity word_replacer_sv_unit is
end word_replacer_sv_unit;
