library verilog;
use verilog.vl_types.all;
entity signextend_sv_unit is
end signextend_sv_unit;
