library verilog;
use verilog.vl_types.all;
entity MP3_tb is
end MP3_tb;
