library verilog;
use verilog.vl_types.all;
entity data_selector_sv_unit is
end data_selector_sv_unit;
