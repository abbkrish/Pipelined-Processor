library verilog;
use verilog.vl_types.all;
entity EX_MEM_register_sv_unit is
end EX_MEM_register_sv_unit;
