library verilog;
use verilog.vl_types.all;
entity zeroextShift_sv_unit is
end zeroextShift_sv_unit;
