library verilog;
use verilog.vl_types.all;
entity cache_hierarchy_sv_unit is
end cache_hierarchy_sv_unit;
