library verilog;
use verilog.vl_types.all;
entity MEM_MEMWB_register_sv_unit is
end MEM_MEMWB_register_sv_unit;
