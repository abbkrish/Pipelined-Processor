library verilog;
use verilog.vl_types.all;
entity addr_splitter_sv_unit is
end addr_splitter_sv_unit;
