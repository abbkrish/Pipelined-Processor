library verilog;
use verilog.vl_types.all;
entity icache_control_sv_unit is
end icache_control_sv_unit;
