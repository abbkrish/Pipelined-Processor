library verilog;
use verilog.vl_types.all;
entity pipeline_datapath_sv_unit is
end pipeline_datapath_sv_unit;
