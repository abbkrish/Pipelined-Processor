library verilog;
use verilog.vl_types.all;
entity shift_sv_unit is
end shift_sv_unit;
