library verilog;
use verilog.vl_types.all;
entity branchAdder_sv_unit is
end branchAdder_sv_unit;
